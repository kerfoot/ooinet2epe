netcdf GP05MOAS-Glider-001-ggldr_dosta_delayed-b373b93231c24b64ac9d79a11bc47078 {
dimensions:
	row = 78737 ;
	preferred_timestamp_strlen = 18 ;
variables:
	double driver_timestamp(row) ;
		driver_timestamp:actual_range = 1391560823.75671, 1394226501.15999 ;
		driver_timestamp:display_name = "Driver Timestamp, seconds since 1900-01-01" ;
		driver_timestamp:internal_name = "driver_timestamp" ;
		driver_timestamp:ioos_category = "Time" ;
		driver_timestamp:long_name = "Driver Timestamp, seconds since 1900-01-01" ;
		driver_timestamp:time_origin = "01-JAN-1970 00:00:00" ;
		driver_timestamp:time_precision = "1970-01-01T00:00:00.000Z" ;
		driver_timestamp:units = "seconds since 1970-01-01T00:00:00Z" ;
	double ingestion_timestamp(row) ;
		ingestion_timestamp:actual_range = 1391560832.13853, 1394226507.67042 ;
		ingestion_timestamp:display_name = "Ingestion Timestamp, seconds since 1900-01-01" ;
		ingestion_timestamp:internal_name = "ingestion_timestamp" ;
		ingestion_timestamp:ioos_category = "Time" ;
		ingestion_timestamp:long_name = "Ingestion Timestamp, seconds since 1900-01-01" ;
		ingestion_timestamp:time_origin = "01-JAN-1970 00:00:00" ;
		ingestion_timestamp:time_precision = "1970-01-01T00:00:00.000Z" ;
		ingestion_timestamp:units = "seconds since 1970-01-01T00:00:00Z" ;
	double internal_timestamp(row) ;
		internal_timestamp:actual_range = 1374259006.3248, 1394193742.25864 ;
		internal_timestamp:display_name = "Internal Timestamp, seconds since 1900-01-01" ;
		internal_timestamp:internal_name = "internal_timestamp" ;
		internal_timestamp:ioos_category = "Time" ;
		internal_timestamp:long_name = "Internal Timestamp, seconds since 1900-01-01" ;
		internal_timestamp:time_origin = "01-JAN-1970 00:00:00" ;
		internal_timestamp:time_precision = "1970-01-01T00:00:00.000Z" ;
		internal_timestamp:units = "seconds since 1970-01-01T00:00:00Z" ;
	float m_present_secs_into_mission(row) ;
		m_present_secs_into_mission:actual_range = 6.21555f, 3160580.f ;
		m_present_secs_into_mission:display_name = "Elapsed mission time, Secs" ;
		m_present_secs_into_mission:internal_name = "m_present_secs_into_mission" ;
		m_present_secs_into_mission:ioos_category = "Dissolved Nutrients" ;
		m_present_secs_into_mission:long_name = "Elapsed mission time, Secs" ;
		m_present_secs_into_mission:precision = "4" ;
		m_present_secs_into_mission:reference_urls = "Gliders" ;
		m_present_secs_into_mission:units = "s" ;
	double m_present_time(row) ;
		m_present_time:actual_range = 1374259006.3248, 1394193742.25864 ;
		m_present_time:display_name = "Time at the start of the cycle, Secs" ;
		m_present_time:internal_name = "m_present_time" ;
		m_present_time:ioos_category = "Time" ;
		m_present_time:long_name = "Time at the start of the cycle, Secs" ;
		m_present_time:precision = "4" ;
		m_present_time:reference_urls = "Gliders" ;
		m_present_time:time_origin = "01-JAN-1970 00:00:00" ;
		m_present_time:time_precision = "1970-01-01T00:00:00.000Z" ;
		m_present_time:units = "seconds since 1970-01-01T00:00:00Z" ;
	char preferred_timestamp(row, preferred_timestamp_strlen) ;
		preferred_timestamp:display_name = "Preferred Timestamp" ;
		preferred_timestamp:internal_name = "preferred_timestamp" ;
		preferred_timestamp:ioos_category = "Time" ;
		preferred_timestamp:long_name = "Preferred Timestamp" ;
		preferred_timestamp:precision = "0" ;
		preferred_timestamp:units = "1" ;
	float sci_m_present_secs_into_mission(row) ;
		sci_m_present_secs_into_mission:actual_range = 6.21555f, 3160580.f ;
		sci_m_present_secs_into_mission:display_name = "Elapsed mission time based on science derived start time, Secs" ;
		sci_m_present_secs_into_mission:internal_name = "sci_m_present_secs_into_mission" ;
		sci_m_present_secs_into_mission:ioos_category = "Dissolved Nutrients" ;
		sci_m_present_secs_into_mission:long_name = "Elapsed mission time based on science derived start time, Secs" ;
		sci_m_present_secs_into_mission:precision = "4" ;
		sci_m_present_secs_into_mission:reference_urls = "Gliders" ;
		sci_m_present_secs_into_mission:units = "s" ;
	double sci_m_present_time(row) ;
		sci_m_present_time:actual_range = 1374259006.3248, 1394193742.25864 ;
		sci_m_present_time:display_name = "Science derived time at the start of the cycle, Secs" ;
		sci_m_present_time:internal_name = "sci_m_present_time" ;
		sci_m_present_time:ioos_category = "Time" ;
		sci_m_present_time:long_name = "Science derived time at the start of the cycle, Secs" ;
		sci_m_present_time:precision = "4" ;
		sci_m_present_time:reference_urls = "Gliders" ;
		sci_m_present_time:time_origin = "01-JAN-1970 00:00:00" ;
		sci_m_present_time:time_precision = "1970-01-01T00:00:00.000Z" ;
		sci_m_present_time:units = "seconds since 1970-01-01T00:00:00Z" ;
	float sci_oxy4_oxygen(row) ;
		sci_oxy4_oxygen:actual_range = 0.f, 304.142f ;
		sci_oxy4_oxygen:display_name = "Estimated Oxygen Concentration, uMol" ;
		sci_oxy4_oxygen:internal_name = "sci_oxy4_oxygen" ;
		sci_oxy4_oxygen:ioos_category = "Dissolved O2" ;
		sci_oxy4_oxygen:long_name = "Estimated Oxygen Concentration, uMol" ;
		sci_oxy4_oxygen:ooi_short_name = "DOCONCS_L1" ;
		sci_oxy4_oxygen:precision = "4" ;
		sci_oxy4_oxygen:reference_urls = "Gliders" ;
		sci_oxy4_oxygen:units = "umol L-1" ;
	float sci_oxy4_saturation(row) ;
		sci_oxy4_saturation:actual_range = 0.f, 105.781f ;
		sci_oxy4_saturation:display_name = "Estimated Percentage Oxygen Saturation, %" ;
		sci_oxy4_saturation:internal_name = "sci_oxy4_saturation" ;
		sci_oxy4_saturation:ioos_category = "Location" ;
		sci_oxy4_saturation:long_name = "Estimated Percentage Oxygen Saturation, %" ;
		sci_oxy4_saturation:precision = "4" ;
		sci_oxy4_saturation:reference_urls = "Gliders" ;
		sci_oxy4_saturation:units = "%" ;
	double time(row) ;
		time:_CoordinateAxisType = "Time" ;
		time:actual_range = 1374259006.3248, 1394193742.25864 ;
		time:axis = "T" ;
		time:display_name = "Time, seconds since 1900-01-01" ;
		time:internal_name = "time" ;
		time:ioos_category = "Time" ;
		time:long_name = "Time, seconds since 1900-01-01" ;
		time:standard_name = "time" ;
		time:time_origin = "01-JAN-1970 00:00:00" ;
		time:time_precision = "1970-01-01T00:00:00.000Z" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;

// global attributes:
		:cdm_data_type = "Other" ;
		:Conventions = "COARDS, CF-1.6, Unidata Dataset Discovery v1.0" ;
		:history = "2014-03-17T18:50:56Z http://sg.b.oceanobservatories.org:10999/5066b4479c4b43279c81c6bd05abf0a5\n",
			"2014-03-17T18:50:56Z http://r2-erddap-prod.oceanobservatories.org:8080/erddap/tabledap/datab373b93231c24b64ac9d79a11bc47078.nc" ;
		:id = "datab373b93231c24b64ac9d79a11bc47078_8571_f367_229e" ;
		:infoUrl = "http://ion-beta.oceanobservatories.org/DataProduct/face/b373b93231c24b64ac9d79a11bc47078" ;
		:institution = "OOI" ;
		:license = "These data were collected by the Ocean Observatory Initiative (OOI) project purely for internal system development purposes during the construction phase of the project and are offered for release to the public with no assurance of data quality, consistency, temporal continuity or additional support. The OOI Program assumes no liability resulting from the use of these data for other than the intended purpose. No data quality assurance steps have been implemented on this data to date." ;
		:sourceUrl = "http://sg.b.oceanobservatories.org:10999/5066b4479c4b43279c81c6bd05abf0a5" ;
		:standard_name_vocabulary = "CF-12" ;
		:summary = "5066b4479c4b43279c81c6bd05abf0a5" ;
		:time_coverage_end = "2014-03-07T12:02:22Z" ;
		:time_coverage_start = "2013-07-19T18:36:46Z" ;
		:title = "Instrument GP05MOAS-GL001-02-DOSTAM999 stream \'ggldr_dosta_delayed\' data product" ;
}
