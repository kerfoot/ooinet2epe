netcdf GP05MOAS-Glider-001-ggldr_eng_delayed-47ae6b72ba644a439a992de4d40c4330 {
dimensions:
	row = 125165 ;
	preferred_timestamp_strlen = 18 ;
variables:
	float c_battpos(row) ;
		c_battpos:actual_range = -9999999.f, 0.7f ;
		c_battpos:display_name = "Commanded Battery Position, inches" ;
		c_battpos:internal_name = "c_battpos" ;
		c_battpos:ioos_category = "Unknown" ;
		c_battpos:long_name = "Commanded Battery Position, inches" ;
		c_battpos:precision = "4" ;
		c_battpos:reference_urls = "Gliders" ;
		c_battpos:units = "in" ;
	float c_wpt_lat(row) ;
		c_wpt_lat:actual_range = -9999999.f, 50.42f ;
		c_wpt_lat:display_name = "Commanded Waypoint Position: Latitude, degrees" ;
		c_wpt_lat:internal_name = "c_wpt_lat" ;
		c_wpt_lat:ioos_category = "Location" ;
		c_wpt_lat:long_name = "Commanded Waypoint Position: Latitude, degrees" ;
		c_wpt_lat:precision = "4" ;
		c_wpt_lat:reference_urls = "Gliders" ;
		c_wpt_lat:units = "degrees" ;
	float c_wpt_lon(row) ;
		c_wpt_lon:actual_range = -9999999.f, -70.53497f ;
		c_wpt_lon:display_name = "Commanded Waypoint Position: Longitude, degrees" ;
		c_wpt_lon:internal_name = "c_wpt_lon" ;
		c_wpt_lon:ioos_category = "Location" ;
		c_wpt_lon:long_name = "Commanded Waypoint Position: Longitude, degrees" ;
		c_wpt_lon:precision = "4" ;
		c_wpt_lon:reference_urls = "Gliders" ;
		c_wpt_lon:units = "degrees" ;
	double driver_timestamp(row) ;
		driver_timestamp:actual_range = 1391560817.66637, 1394226503.41514 ;
		driver_timestamp:display_name = "Driver Timestamp, seconds since 1900-01-01" ;
		driver_timestamp:internal_name = "driver_timestamp" ;
		driver_timestamp:ioos_category = "Time" ;
		driver_timestamp:long_name = "Driver Timestamp, seconds since 1900-01-01" ;
		driver_timestamp:time_origin = "01-JAN-1970 00:00:00" ;
		driver_timestamp:time_precision = "1970-01-01T00:00:00.000Z" ;
		driver_timestamp:units = "seconds since 1970-01-01T00:00:00Z" ;
	double ingestion_timestamp(row) ;
		ingestion_timestamp:actual_range = 1391560827.00056, 1394226517.27003 ;
		ingestion_timestamp:display_name = "Ingestion Timestamp, seconds since 1900-01-01" ;
		ingestion_timestamp:internal_name = "ingestion_timestamp" ;
		ingestion_timestamp:ioos_category = "Time" ;
		ingestion_timestamp:long_name = "Ingestion Timestamp, seconds since 1900-01-01" ;
		ingestion_timestamp:time_origin = "01-JAN-1970 00:00:00" ;
		ingestion_timestamp:time_precision = "1970-01-01T00:00:00.000Z" ;
		ingestion_timestamp:units = "seconds since 1970-01-01T00:00:00Z" ;
	double internal_timestamp(row) ;
		internal_timestamp:actual_range = 1374259009.34088, 1394223427.29788 ;
		internal_timestamp:display_name = "Internal Timestamp, seconds since 1900-01-01" ;
		internal_timestamp:internal_name = "internal_timestamp" ;
		internal_timestamp:ioos_category = "Time" ;
		internal_timestamp:long_name = "Internal Timestamp, seconds since 1900-01-01" ;
		internal_timestamp:time_origin = "01-JAN-1970 00:00:00" ;
		internal_timestamp:time_precision = "1970-01-01T00:00:00.000Z" ;
		internal_timestamp:units = "seconds since 1970-01-01T00:00:00Z" ;
	float m_battpos(row) ;
		m_battpos:actual_range = -9999999.f, 0.725462f ;
		m_battpos:display_name = "Measured Battery Position, inches" ;
		m_battpos:internal_name = "m_battpos" ;
		m_battpos:ioos_category = "Unknown" ;
		m_battpos:long_name = "Measured Battery Position, inches" ;
		m_battpos:precision = "4" ;
		m_battpos:reference_urls = "Gliders" ;
		m_battpos:units = "in" ;
	float m_coulomb_amphr_total(row) ;
		m_coulomb_amphr_total:actual_range = -9999999.f, 673.741f ;
		m_coulomb_amphr_total:display_name = "Measured Total Persistant amp-hours, Ah" ;
		m_coulomb_amphr_total:internal_name = "m_coulomb_amphr_total" ;
		m_coulomb_amphr_total:ioos_category = "Salinity" ;
		m_coulomb_amphr_total:long_name = "Measured Total Persistant amp-hours, Ah" ;
		m_coulomb_amphr_total:precision = "4" ;
		m_coulomb_amphr_total:reference_urls = "Gliders" ;
		m_coulomb_amphr_total:units = "amp-h" ;
	float m_coulomb_current(row) ;
		m_coulomb_current:actual_range = -9999999.f, 5.84517f ;
		m_coulomb_current:display_name = "Measured Instantaneous Current, A" ;
		m_coulomb_current:internal_name = "m_coulomb_current" ;
		m_coulomb_current:ioos_category = "Currents" ;
		m_coulomb_current:long_name = "Measured Instantaneous Current, A" ;
		m_coulomb_current:precision = "4" ;
		m_coulomb_current:reference_urls = "Gliders" ;
		m_coulomb_current:units = "amp" ;
	float m_de_oil_vol(row) ;
		m_de_oil_vol:actual_range = -9999999.f, 261.613f ;
		m_de_oil_vol:display_name = "Measured Deep Electric Oil Volume, mL" ;
		m_de_oil_vol:internal_name = "m_de_oil_vol" ;
		m_de_oil_vol:ioos_category = "Unknown" ;
		m_de_oil_vol:long_name = "Measured Deep Electric Oil Volume, mL" ;
		m_de_oil_vol:precision = "4" ;
		m_de_oil_vol:reference_urls = "Gliders" ;
		m_de_oil_vol:units = "mL" ;
	float m_depth(row) ;
		m_depth:actual_range = -9999999.f, 978.424f ;
		m_depth:display_name = "Measured Depth, m" ;
		m_depth:internal_name = "m_depth" ;
		m_depth:ioos_category = "Location" ;
		m_depth:long_name = "Measured Depth, m" ;
		m_depth:precision = "4" ;
		m_depth:reference_urls = "Gliders" ;
		m_depth:units = "m" ;
	float m_gps_lat(row) ;
		m_gps_lat:actual_range = -9999999.f, 2312.15f ;
		m_gps_lat:display_name = "Measured GPS Latitude, degrees" ;
		m_gps_lat:internal_name = "m_gps_lat" ;
		m_gps_lat:ioos_category = "Location" ;
		m_gps_lat:long_name = "Measured GPS Latitude, degrees" ;
		m_gps_lat:precision = "4" ;
		m_gps_lat:reference_urls = "Gliders" ;
		m_gps_lat:units = "degrees" ;
	float m_gps_lon(row) ;
		m_gps_lon:actual_range = -9999999.f, 2312.15f ;
		m_gps_lon:display_name = "Measured GPS Longitude, degrees" ;
		m_gps_lon:internal_name = "m_gps_lon" ;
		m_gps_lon:ioos_category = "Location" ;
		m_gps_lon:long_name = "Measured GPS Longitude, degrees" ;
		m_gps_lon:precision = "4" ;
		m_gps_lon:reference_urls = "Gliders" ;
		m_gps_lon:units = "degrees" ;
	float m_heading(row) ;
		m_heading:actual_range = -9999999.f, 6.28144f ;
		m_heading:display_name = "Measured Heading, rad" ;
		m_heading:internal_name = "m_heading" ;
		m_heading:ioos_category = "Unknown" ;
		m_heading:long_name = "Measured Heading, rad" ;
		m_heading:precision = "4" ;
		m_heading:reference_urls = "Gliders" ;
		m_heading:units = "rad" ;
	float m_lat(row) ;
		m_lat:actual_range = -9999999.f, 50.90302f ;
		m_lat:display_name = "Derived latitude, degrees" ;
		m_lat:internal_name = "m_lat" ;
		m_lat:ioos_category = "Location" ;
		m_lat:long_name = "Derived latitude, degrees" ;
		m_lat:precision = "4" ;
		m_lat:reference_urls = "Gliders" ;
		m_lat:units = "degrees" ;
	float m_lon(row) ;
		m_lon:actual_range = -9999999.f, -70.53497f ;
		m_lon:display_name = "Derived longitude, degrees" ;
		m_lon:internal_name = "m_lon" ;
		m_lon:ioos_category = "Location" ;
		m_lon:long_name = "Derived longitude, degrees" ;
		m_lon:precision = "4" ;
		m_lon:reference_urls = "Gliders" ;
		m_lon:units = "degrees" ;
	float m_pitch(row) ;
		m_pitch:actual_range = -9999999.f, 1.03149f ;
		m_pitch:display_name = "Measured Pitch, Radians" ;
		m_pitch:internal_name = "m_pitch" ;
		m_pitch:ioos_category = "Identifier" ;
		m_pitch:long_name = "Measured Pitch, Radians" ;
		m_pitch:precision = "4" ;
		m_pitch:reference_urls = "Gliders" ;
		m_pitch:units = "rad" ;
	float m_present_secs_into_mission(row) ;
		m_present_secs_into_mission:actual_range = 0.f, 3190230.f ;
		m_present_secs_into_mission:display_name = "Elapsed mission time, Secs" ;
		m_present_secs_into_mission:internal_name = "m_present_secs_into_mission" ;
		m_present_secs_into_mission:ioos_category = "Dissolved Nutrients" ;
		m_present_secs_into_mission:long_name = "Elapsed mission time, Secs" ;
		m_present_secs_into_mission:precision = "4" ;
		m_present_secs_into_mission:reference_urls = "Gliders" ;
		m_present_secs_into_mission:units = "s" ;
	double m_present_time(row) ;
		m_present_time:actual_range = 1374259009.34088, 1394223427.29788 ;
		m_present_time:display_name = "Time at the start of the cycle, Secs" ;
		m_present_time:internal_name = "m_present_time" ;
		m_present_time:ioos_category = "Time" ;
		m_present_time:long_name = "Time at the start of the cycle, Secs" ;
		m_present_time:precision = "4" ;
		m_present_time:reference_urls = "Gliders" ;
		m_present_time:time_origin = "01-JAN-1970 00:00:00" ;
		m_present_time:time_precision = "1970-01-01T00:00:00.000Z" ;
		m_present_time:units = "seconds since 1970-01-01T00:00:00Z" ;
	float m_speed(row) ;
		m_speed:actual_range = -9999999.f, 0.537062f ;
		m_speed:display_name = "Measured Speed, m/s" ;
		m_speed:internal_name = "m_speed" ;
		m_speed:ioos_category = "Unknown" ;
		m_speed:long_name = "Measured Speed, m/s" ;
		m_speed:precision = "4" ;
		m_speed:reference_urls = "Gliders" ;
		m_speed:units = "m s-1" ;
	float m_water_vx(row) ;
		m_water_vx:actual_range = -9999999.f, 2.04297f ;
		m_water_vx:display_name = "Measured Water Velocity: X, m/s" ;
		m_water_vx:internal_name = "m_water_vx" ;
		m_water_vx:ioos_category = "Location" ;
		m_water_vx:long_name = "Measured Water Velocity: X, m/s" ;
		m_water_vx:precision = "4" ;
		m_water_vx:reference_urls = "Gliders" ;
		m_water_vx:units = "m s-1" ;
	float m_water_vy(row) ;
		m_water_vy:actual_range = -9999999.f, 2.65241f ;
		m_water_vy:display_name = "Measured Water Velocity: Y, m/s" ;
		m_water_vy:internal_name = "m_water_vy" ;
		m_water_vy:ioos_category = "Location" ;
		m_water_vy:long_name = "Measured Water Velocity: Y, m/s" ;
		m_water_vy:precision = "4" ;
		m_water_vy:reference_urls = "Gliders" ;
		m_water_vy:units = "m s-1" ;
	char preferred_timestamp(row, preferred_timestamp_strlen) ;
		preferred_timestamp:display_name = "Preferred Timestamp" ;
		preferred_timestamp:internal_name = "preferred_timestamp" ;
		preferred_timestamp:ioos_category = "Time" ;
		preferred_timestamp:long_name = "Preferred Timestamp" ;
		preferred_timestamp:precision = "0" ;
		preferred_timestamp:units = "1" ;
	double time(row) ;
		time:_CoordinateAxisType = "Time" ;
		time:actual_range = 1374259009.34088, 1394223427.29788 ;
		time:axis = "T" ;
		time:display_name = "Time, seconds since 1900-01-01" ;
		time:internal_name = "time" ;
		time:ioos_category = "Time" ;
		time:long_name = "Time, seconds since 1900-01-01" ;
		time:standard_name = "time" ;
		time:time_origin = "01-JAN-1970 00:00:00" ;
		time:time_precision = "1970-01-01T00:00:00.000Z" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
	float x_low_power_status(row) ;
		x_low_power_status:actual_range = -9999999.f, 13.f ;
		x_low_power_status:display_name = "Low Power Status" ;
		x_low_power_status:internal_name = "x_low_power_status" ;
		x_low_power_status:ioos_category = "Location" ;
		x_low_power_status:long_name = "Low Power Status" ;
		x_low_power_status:precision = "4" ;
		x_low_power_status:reference_urls = "Gliders" ;
		x_low_power_status:units = "1" ;

// global attributes:
		:cdm_data_type = "Other" ;
		:Conventions = "COARDS, CF-1.6, Unidata Dataset Discovery v1.0" ;
		:history = "2014-03-17T18:51:51Z http://sg.b.oceanobservatories.org:10999/3db0d8e176af4ce384da7bffd3334ab0\n",
			"2014-03-17T18:51:51Z http://r2-erddap-prod.oceanobservatories.org:8080/erddap/tabledap/data47ae6b72ba644a439a992de4d40c4330.nc" ;
		:id = "data47ae6b72ba644a439a992de4d40c4330_8571_f367_229e" ;
		:infoUrl = "http://ion-beta.oceanobservatories.org/DataProduct/face/47ae6b72ba644a439a992de4d40c4330" ;
		:institution = "OOI" ;
		:license = "These data were collected by the Ocean Observatory Initiative (OOI) project purely for internal system development purposes during the construction phase of the project and are offered for release to the public with no assurance of data quality, consistency, temporal continuity or additional support. The OOI Program assumes no liability resulting from the use of these data for other than the intended purpose. No data quality assurance steps have been implemented on this data to date." ;
		:sourceUrl = "http://sg.b.oceanobservatories.org:10999/3db0d8e176af4ce384da7bffd3334ab0" ;
		:standard_name_vocabulary = "CF-12" ;
		:summary = "3db0d8e176af4ce384da7bffd3334ab0" ;
		:time_coverage_end = "2014-03-07T20:17:07Z" ;
		:time_coverage_start = "2013-07-19T18:36:49Z" ;
		:title = "Platform GP05MOAS-GL001 stream \'ggldr_eng_delayed\' data product" ;
}
