netcdf GP05MOAS-Glider-001-FLUBSCT-44e6943f323f4938b78311f49593f66d {
dimensions:
	row = 74241 ;
variables:
	float sci_flbb_bb_units(row) ;
		sci_flbb_bb_units:actual_range = 0.f, 0.0057113f ;
		sci_flbb_bb_units:display_name = "Volume Scattering Function, Beta(117,650), m-1 sr-1" ;
		sci_flbb_bb_units:internal_name = "sci_flbb_bb_units" ;
		sci_flbb_bb_units:ioos_category = "Unknown" ;
		sci_flbb_bb_units:long_name = "Volume Scattering Function, Beta(117,650), m-1 sr-1" ;
		sci_flbb_bb_units:ooi_short_name = "FLUBSCT_L1" ;
		sci_flbb_bb_units:precision = "4" ;
		sci_flbb_bb_units:reference_urls = "Gliders" ;
		sci_flbb_bb_units:units = "m-1 sr-1" ;
	double time(row) ;
		time:_CoordinateAxisType = "Time" ;
		time:actual_range = 1374259006.3248, 1394193738.24521 ;
		time:axis = "T" ;
		time:display_name = "Time, seconds since 1900-01-01" ;
		time:internal_name = "time" ;
		time:ioos_category = "Time" ;
		time:long_name = "Time, seconds since 1900-01-01" ;
		time:standard_name = "time" ;
		time:time_origin = "01-JAN-1970 00:00:00" ;
		time:time_precision = "1970-01-01T00:00:00.000Z" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;

// global attributes:
		:cdm_data_type = "Other" ;
		:Conventions = "COARDS, CF-1.6, Unidata Dataset Discovery v1.0" ;
		:history = "2014-03-17T18:51:59Z http://sg.b.oceanobservatories.org:10999/86f942d089b749c7b630304f4cf212ad\n",
			"2014-03-17T18:51:59Z http://r2-erddap-prod.oceanobservatories.org:8080/erddap/tabledap/data44e6943f323f4938b78311f49593f66d.nc" ;
		:id = "data44e6943f323f4938b78311f49593f66d_8571_f367_229e" ;
		:infoUrl = "http://ion-beta.oceanobservatories.org/DataProduct/face/44e6943f323f4938b78311f49593f66d" ;
		:institution = "OOI" ;
		:license = "These data were collected by the Ocean Observatory Initiative (OOI) project purely for internal system development purposes during the construction phase of the project and are offered for release to the public with no assurance of data quality, consistency, temporal continuity or additional support. The OOI Program assumes no liability resulting from the use of these data for other than the intended purpose. No data quality assurance steps have been implemented on this data to date." ;
		:sourceUrl = "http://sg.b.oceanobservatories.org:10999/86f942d089b749c7b630304f4cf212ad" ;
		:standard_name_vocabulary = "CF-12" ;
		:summary = "86f942d089b749c7b630304f4cf212ad" ;
		:time_coverage_end = "2014-03-07T12:02:18Z" ;
		:time_coverage_start = "2013-07-19T18:36:46Z" ;
		:title = "Optical Backscatter (Red Wavelengths) L1 FLORD Glider 001 - Global Station Papa Mobile Assets" ;
}
