netcdf GP05MOAS-Glider-001-ggldr_ctdgv_delayed-0b9b23e7ae8c495bb6f6f36fc29b1ec0 {
dimensions:
	row = 78719 ;
	preferred_timestamp_strlen = 18 ;
variables:
	byte cmbnflg_qc(row) ;
		cmbnflg_qc:actual_range = 0b, 0b ;
		cmbnflg_qc:display_name = "Combined Data Quality Control Flag" ;
		cmbnflg_qc:ioos_category = "Quality" ;
		cmbnflg_qc:long_name = "Combined Data Quality Control Flag" ;
		cmbnflg_qc:ooi_short_name = "CMBNFLG_QC" ;
		cmbnflg_qc:units = "1" ;
	double driver_timestamp(row) ;
		driver_timestamp:actual_range = 1391560835.10617, 1394226500.28635 ;
		driver_timestamp:display_name = "Driver Timestamp, seconds since 1900-01-01" ;
		driver_timestamp:internal_name = "driver_timestamp" ;
		driver_timestamp:ioos_category = "Time" ;
		driver_timestamp:long_name = "Driver Timestamp, seconds since 1900-01-01" ;
		driver_timestamp:time_origin = "01-JAN-1970 00:00:00" ;
		driver_timestamp:time_precision = "1970-01-01T00:00:00.000Z" ;
		driver_timestamp:units = "seconds since 1970-01-01T00:00:00Z" ;
	double ingestion_timestamp(row) ;
		ingestion_timestamp:actual_range = 1391560844.55446, 1394226513.79987 ;
		ingestion_timestamp:display_name = "Ingestion Timestamp, seconds since 1900-01-01" ;
		ingestion_timestamp:internal_name = "ingestion_timestamp" ;
		ingestion_timestamp:ioos_category = "Time" ;
		ingestion_timestamp:long_name = "Ingestion Timestamp, seconds since 1900-01-01" ;
		ingestion_timestamp:time_origin = "01-JAN-1970 00:00:00" ;
		ingestion_timestamp:time_precision = "1970-01-01T00:00:00.000Z" ;
		ingestion_timestamp:units = "seconds since 1970-01-01T00:00:00Z" ;
	double internal_timestamp(row) ;
		internal_timestamp:actual_range = 1374259006.3248, 1394193745.27017 ;
		internal_timestamp:display_name = "Internal Timestamp, seconds since 1900-01-01" ;
		internal_timestamp:internal_name = "internal_timestamp" ;
		internal_timestamp:ioos_category = "Time" ;
		internal_timestamp:long_name = "Internal Timestamp, seconds since 1900-01-01" ;
		internal_timestamp:time_origin = "01-JAN-1970 00:00:00" ;
		internal_timestamp:time_precision = "1970-01-01T00:00:00.000Z" ;
		internal_timestamp:units = "seconds since 1970-01-01T00:00:00Z" ;
	float m_present_secs_into_mission(row) ;
		m_present_secs_into_mission:actual_range = 6.21555f, 3160580.f ;
		m_present_secs_into_mission:display_name = "Elapsed mission time, Secs" ;
		m_present_secs_into_mission:internal_name = "m_present_secs_into_mission" ;
		m_present_secs_into_mission:ioos_category = "Dissolved Nutrients" ;
		m_present_secs_into_mission:long_name = "Elapsed mission time, Secs" ;
		m_present_secs_into_mission:precision = "4" ;
		m_present_secs_into_mission:reference_urls = "Gliders" ;
		m_present_secs_into_mission:units = "s" ;
	double m_present_time(row) ;
		m_present_time:actual_range = 1374259006.3248, 1394193745.27017 ;
		m_present_time:display_name = "Time at the start of the cycle, Secs" ;
		m_present_time:internal_name = "m_present_time" ;
		m_present_time:ioos_category = "Time" ;
		m_present_time:long_name = "Time at the start of the cycle, Secs" ;
		m_present_time:precision = "4" ;
		m_present_time:reference_urls = "Gliders" ;
		m_present_time:time_origin = "01-JAN-1970 00:00:00" ;
		m_present_time:time_precision = "1970-01-01T00:00:00.000Z" ;
		m_present_time:units = "seconds since 1970-01-01T00:00:00Z" ;
	byte pracsal_glblrng_qc(row) ;
		pracsal_glblrng_qc:actual_range = 0b, 0b ;
		pracsal_glblrng_qc:display_name = "PRACSAL Global Range Test Quality Control Flag" ;
		pracsal_glblrng_qc:ioos_category = "Quality" ;
		pracsal_glblrng_qc:long_name = "PRACSAL Global Range Test Quality Control Flag" ;
		pracsal_glblrng_qc:ooi_short_name = "PRACSAL_GLBLRNG_QC" ;
		pracsal_glblrng_qc:units = "1" ;
	byte pracsal_gradtst_qc(row) ;
		pracsal_gradtst_qc:actual_range = 0b, 0b ;
		pracsal_gradtst_qc:display_name = "PRACSAL Gradient Test Quality Control Flag" ;
		pracsal_gradtst_qc:ioos_category = "Quality" ;
		pracsal_gradtst_qc:long_name = "PRACSAL Gradient Test Quality Control Flag" ;
		pracsal_gradtst_qc:ooi_short_name = "PRACSAL_GRADTST_QC" ;
		pracsal_gradtst_qc:units = "1" ;
	byte pracsal_loclrng_qc(row) ;
		pracsal_loclrng_qc:actual_range = 0b, 0b ;
		pracsal_loclrng_qc:display_name = "PRACSAL Local Range Test Quality Control Flag" ;
		pracsal_loclrng_qc:ioos_category = "Quality" ;
		pracsal_loclrng_qc:long_name = "PRACSAL Local Range Test Quality Control Flag" ;
		pracsal_loclrng_qc:ooi_short_name = "PRACSAL_LOCLRNG_QC" ;
		pracsal_loclrng_qc:units = "1" ;
	byte pracsal_spketst_qc(row) ;
		pracsal_spketst_qc:actual_range = 0b, 0b ;
		pracsal_spketst_qc:display_name = "PRACSAL Spike Test Quality Control Flag" ;
		pracsal_spketst_qc:ioos_category = "Quality" ;
		pracsal_spketst_qc:long_name = "PRACSAL Spike Test Quality Control Flag" ;
		pracsal_spketst_qc:ooi_short_name = "PRACSAL_SPKETST_QC" ;
		pracsal_spketst_qc:units = "1" ;
	byte pracsal_stuckvl_qc(row) ;
		pracsal_stuckvl_qc:actual_range = 0b, 0b ;
		pracsal_stuckvl_qc:display_name = "PRACSAL Stuck Value Test Quality Control Flag" ;
		pracsal_stuckvl_qc:ioos_category = "Quality" ;
		pracsal_stuckvl_qc:long_name = "PRACSAL Stuck Value Test Quality Control Flag" ;
		pracsal_stuckvl_qc:ooi_short_name = "PRACSAL_STUCKVL_QC" ;
		pracsal_stuckvl_qc:units = "1" ;
	char preferred_timestamp(row, preferred_timestamp_strlen) ;
		preferred_timestamp:display_name = "Preferred Timestamp" ;
		preferred_timestamp:internal_name = "preferred_timestamp" ;
		preferred_timestamp:ioos_category = "Time" ;
		preferred_timestamp:long_name = "Preferred Timestamp" ;
		preferred_timestamp:precision = "0" ;
		preferred_timestamp:units = "1" ;
	float sci_m_present_secs_into_mission(row) ;
		sci_m_present_secs_into_mission:actual_range = 6.21555f, 3160580.f ;
		sci_m_present_secs_into_mission:display_name = "Elapsed mission time based on science derived start time, Secs" ;
		sci_m_present_secs_into_mission:internal_name = "sci_m_present_secs_into_mission" ;
		sci_m_present_secs_into_mission:ioos_category = "Dissolved Nutrients" ;
		sci_m_present_secs_into_mission:long_name = "Elapsed mission time based on science derived start time, Secs" ;
		sci_m_present_secs_into_mission:precision = "4" ;
		sci_m_present_secs_into_mission:reference_urls = "Gliders" ;
		sci_m_present_secs_into_mission:units = "s" ;
	double sci_m_present_time(row) ;
		sci_m_present_time:actual_range = 1374259006.3248, 1394193745.27017 ;
		sci_m_present_time:display_name = "Science derived time at the start of the cycle, Secs" ;
		sci_m_present_time:internal_name = "sci_m_present_time" ;
		sci_m_present_time:ioos_category = "Time" ;
		sci_m_present_time:long_name = "Science derived time at the start of the cycle, Secs" ;
		sci_m_present_time:precision = "4" ;
		sci_m_present_time:reference_urls = "Gliders" ;
		sci_m_present_time:time_origin = "01-JAN-1970 00:00:00" ;
		sci_m_present_time:time_precision = "1970-01-01T00:00:00.000Z" ;
		sci_m_present_time:units = "seconds since 1970-01-01T00:00:00Z" ;
	double sci_water_cond(row) ;
		sci_water_cond:actual_range = 0., 4.09281 ;
		sci_water_cond:display_name = "Conductivity, S/m" ;
		sci_water_cond:internal_name = "sci_water_cond" ;
		sci_water_cond:ioos_category = "Unknown" ;
		sci_water_cond:long_name = "Conductivity, S/m" ;
		sci_water_cond:ooi_short_name = "CONDWAT_L1" ;
		sci_water_cond:precision = "4" ;
		sci_water_cond:reference_urls = "Gliders" ;
		sci_water_cond:units = "S m-1" ;
	float sci_water_pracsal(row) ;
		sci_water_pracsal:actual_range = 0.f, 34.86565f ;
		sci_water_pracsal:display_name = "sci_water_pracsal" ;
		sci_water_pracsal:internal_name = "sci_water_pracsal" ;
		sci_water_pracsal:ioos_category = "Unknown" ;
		sci_water_pracsal:long_name = "sci_water_pracsal" ;
		sci_water_pracsal:ooi_short_name = "PRACSAL_L2" ;
		sci_water_pracsal:precision = "4" ;
		sci_water_pracsal:reference_urls = "Gliders" ;
		sci_water_pracsal:units = "1" ;
	double sci_water_pressure(row) ;
		sci_water_pressure:actual_range = -0.024, 99.37 ;
		sci_water_pressure:display_name = "Pressure, bars" ;
		sci_water_pressure:internal_name = "sci_water_pressure" ;
		sci_water_pressure:ioos_category = "Pressure" ;
		sci_water_pressure:long_name = "Pressure, bars" ;
		sci_water_pressure:ooi_short_name = "PRESWAT_L1" ;
		sci_water_pressure:precision = "4" ;
		sci_water_pressure:reference_urls = "Gliders" ;
		sci_water_pressure:units = "bar" ;
	double sci_water_temp(row) ;
		sci_water_temp:actual_range = 0., 21.3943 ;
		sci_water_temp:display_name = "Temperature, degrees C" ;
		sci_water_temp:internal_name = "sci_water_temp" ;
		sci_water_temp:ioos_category = "Temperature" ;
		sci_water_temp:long_name = "Temperature, degrees C" ;
		sci_water_temp:ooi_short_name = "TEMPWAT_L1" ;
		sci_water_temp:precision = "4" ;
		sci_water_temp:reference_urls = "Gliders" ;
		sci_water_temp:units = "deg_C" ;
	double time(row) ;
		time:_CoordinateAxisType = "Time" ;
		time:actual_range = 1374259006.3248, 1394193745.27017 ;
		time:axis = "T" ;
		time:display_name = "Time, seconds since 1900-01-01" ;
		time:internal_name = "time" ;
		time:ioos_category = "Time" ;
		time:long_name = "Time, seconds since 1900-01-01" ;
		time:standard_name = "time" ;
		time:time_origin = "01-JAN-1970 00:00:00" ;
		time:time_precision = "1970-01-01T00:00:00.000Z" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;

// global attributes:
		:cdm_data_type = "Other" ;
		:Conventions = "COARDS, CF-1.6, Unidata Dataset Discovery v1.0" ;
		:history = "2014-03-17T18:51:19Z http://sg.b.oceanobservatories.org:10999/99acf532886d4fb5aaab151d0975917a\n",
			"2014-03-17T18:51:19Z http://r2-erddap-prod.oceanobservatories.org:8080/erddap/tabledap/data0b9b23e7ae8c495bb6f6f36fc29b1ec0.nc" ;
		:id = "data0b9b23e7ae8c495bb6f6f36fc29b1ec0_8571_f367_229e" ;
		:infoUrl = "http://ion-beta.oceanobservatories.org/DataProduct/face/0b9b23e7ae8c495bb6f6f36fc29b1ec0" ;
		:institution = "OOI" ;
		:license = "These data were collected by the Ocean Observatory Initiative (OOI) project purely for internal system development purposes during the construction phase of the project and are offered for release to the public with no assurance of data quality, consistency, temporal continuity or additional support. The OOI Program assumes no liability resulting from the use of these data for other than the intended purpose. No data quality assurance steps have been implemented on this data to date." ;
		:sourceUrl = "http://sg.b.oceanobservatories.org:10999/99acf532886d4fb5aaab151d0975917a" ;
		:standard_name_vocabulary = "CF-12" ;
		:summary = "99acf532886d4fb5aaab151d0975917a" ;
		:time_coverage_end = "2014-03-07T12:02:25Z" ;
		:time_coverage_start = "2013-07-19T18:36:46Z" ;
		:title = "Instrument GP05MOAS-GL001-04-CTDGVM999 stream \'ggldr_ctdgv_delayed\' data product" ;
}
