netcdf GP05MOAS-Glider-001-DOCONCS-e6bca04956e541128a75c1b2f1664e2a {
dimensions:
	row = 78737 ;
variables:
	float sci_oxy4_oxygen(row) ;
		sci_oxy4_oxygen:actual_range = 0.f, 304.142f ;
		sci_oxy4_oxygen:display_name = "Estimated Oxygen Concentration, uMol" ;
		sci_oxy4_oxygen:internal_name = "sci_oxy4_oxygen" ;
		sci_oxy4_oxygen:ioos_category = "Dissolved O2" ;
		sci_oxy4_oxygen:long_name = "Estimated Oxygen Concentration, uMol" ;
		sci_oxy4_oxygen:ooi_short_name = "DOCONCS_L1" ;
		sci_oxy4_oxygen:precision = "4" ;
		sci_oxy4_oxygen:reference_urls = "Gliders" ;
		sci_oxy4_oxygen:units = "umol L-1" ;
	double time(row) ;
		time:_CoordinateAxisType = "Time" ;
		time:actual_range = 1374259006.3248, 1394193742.25864 ;
		time:axis = "T" ;
		time:display_name = "Time, seconds since 1900-01-01" ;
		time:internal_name = "time" ;
		time:ioos_category = "Time" ;
		time:long_name = "Time, seconds since 1900-01-01" ;
		time:standard_name = "time" ;
		time:time_origin = "01-JAN-1970 00:00:00" ;
		time:time_precision = "1970-01-01T00:00:00.000Z" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;

// global attributes:
		:cdm_data_type = "Other" ;
		:Conventions = "COARDS, CF-1.6, Unidata Dataset Discovery v1.0" ;
		:history = "2014-03-17T18:50:30Z http://sg.b.oceanobservatories.org:10999/5066b4479c4b43279c81c6bd05abf0a5\n",
			"2014-03-17T18:50:30Z http://r2-erddap-prod.oceanobservatories.org:8080/erddap/tabledap/datae6bca04956e541128a75c1b2f1664e2a.nc" ;
		:id = "datae6bca04956e541128a75c1b2f1664e2a_8571_f367_229e" ;
		:infoUrl = "http://ion-beta.oceanobservatories.org/DataProduct/face/e6bca04956e541128a75c1b2f1664e2a" ;
		:institution = "OOI" ;
		:license = "These data were collected by the Ocean Observatory Initiative (OOI) project purely for internal system development purposes during the construction phase of the project and are offered for release to the public with no assurance of data quality, consistency, temporal continuity or additional support. The OOI Program assumes no liability resulting from the use of these data for other than the intended purpose. No data quality assurance steps have been implemented on this data to date." ;
		:sourceUrl = "http://sg.b.oceanobservatories.org:10999/5066b4479c4b43279c81c6bd05abf0a5" ;
		:standard_name_vocabulary = "CF-12" ;
		:summary = "5066b4479c4b43279c81c6bd05abf0a5" ;
		:time_coverage_end = "2014-03-07T12:02:22Z" ;
		:time_coverage_start = "2013-07-19T18:36:46Z" ;
		:title = "Oxygen Concentration from Stable DO Instrument L1 DOSTA Glider 001 - Global Station Papa Mobile Assets" ;
}
