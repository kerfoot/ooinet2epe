netcdf GP05MOAS-GL001-20140307T0953 {
dimensions:
	time = 130 ;
	traj_strlen = 14 ;
variables:
	double time(time) ;
		time:ancillary_variables = "" ;
		time:long_name = "Time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
	char trajectory(traj_strlen) ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:comment = "A trajectory is a glider deployment" ;
		trajectory:long_name = "Trajectory Name" ;
		trajectory:units = "1" ;
	double lat(time) ;
		lat:long_name = "Latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = -999. ;
	double lon(time) ;
		lon:long_name = "Longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = -999. ;
	double pressure(time) ;
		pressure:instrument = "instrument_ctd" ;
		pressure:long_name = "Pressure, dbar" ;
		pressure:observation_type = "calculated" ;
		pressure:positive = "down" ;
		pressure:reference_datum = "sea-surface" ;
		pressure:standard_name = "sea_water_pressure" ;
		pressure:units = "dbar" ;
		pressure:valid_max = 2000. ;
		pressure:valid_min = 0. ;
		pressure:_FillValue = -999. ;
	double depth(time) ;
		depth:comment = "" ;
		depth:instrument = "instrument_ctd" ;
		depth:long_name = "Depth, m" ;
		depth:observation_type = "calculated" ;
		depth:positive = "down" ;
		depth:reference_datum = "sea-surface" ;
		depth:standard_name = "depth" ;
		depth:units = "meters" ;
		depth:valid_max = 2000. ;
		depth:valid_min = 0. ;
		depth:_FillValue = -999. ;
	double temperature(time) ;
		temperature:instrument = "instrument_ctd" ;
		temperature:long_name = "Temperature, Celsius" ;
		temperature:observation_type = "measured" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "Celsius" ;
		temperature:valid_max = 40. ;
		temperature:valid_min = -5. ;
		temperature:_FillValue = -999. ;
	double conductivity(time) ;
		conductivity:instrument = "instrument_ctd" ;
		conductivity:long_name = "Conductivity, S m-1" ;
		conductivity:observation_type = "measured" ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:units = "S m-1" ;
		conductivity:valid_max = 10. ;
		conductivity:valid_min = 0. ;
		conductivity:_FillValue = -999. ;
	double salinity(time) ;
		salinity:instrument = "instrument_ctd" ;
		salinity:long_name = "Salinity, PSU" ;
		salinity:observation_type = "calculated" ;
		salinity:standard_name = "sea_water_salinity" ;
		salinity:units = "1" ;
		salinity:valid_max = 40. ;
		salinity:valid_min = 0. ;
		salinity:_FillValue = -999. ;
	double density(time) ;
		density:instrument = "instrument_ctd" ;
		density:long_name = "Density, kg m-3" ;
		density:observation_type = "calculated" ;
		density:standard_name = "sea_water_density" ;
		density:units = "kg m-3" ;
		density:valid_max = 1040. ;
		density:valid_min = 1015. ;
		density:_FillValue = -999. ;
	double chla(time) ;
		chla:instrument = "instrument_flbb" ;
		chla:long_name = "Chlorophyll a Concentration, ug L-1" ;
		chla:observation_type = "measured" ;
		chla:standard_name = "mass_concentration_of_chlorophyll_a_in_sea_water" ;
		chla:units = "ug L-1" ;
		chla:valid_max = 20. ;
		chla:valid_min = 0. ;
		chla:_FillValue = -999. ;
	double bb(time) ;
		bb:instrument = "instrument_flbb" ;
		bb:long_name = "Volume Scattering Function, Beta(117,650), m-1 sr-1" ;
		bb:observation_type = "measured" ;
		bb:units = "m-1 sr-1" ;
		bb:valid_max = 0.1 ;
		bb:valid_min = 0. ;
		bb:_FillValue = -999. ;
	double oxygen_sat(time) ;
		oxygen_sat:instrument = "instrument_optode" ;
		oxygen_sat:long_name = "Estimated Percentage Oxygen Saturation, %" ;
		oxygen_sat:observation_type = "measured" ;
		oxygen_sat:standard_name = "fractional_saturation_of_oxygen_in_sea_water" ;
		oxygen_sat:units = "%" ;
		oxygen_sat:valid_max = 120. ;
		oxygen_sat:valid_min = 0. ;
		oxygen_sat:_FillValue = -999. ;
	double oxygen_conc(time) ;
		oxygen_conc:instrument = "instrument_optode" ;
		oxygen_conc:long_name = "Estimated Oxygen Concentration, uMol L-1" ;
		oxygen_conc:observation_type = "measured" ;
		oxygen_conc:standard_name = "mole_concentration_of_dissolved_molecular_oxygen_in_sea_water" ;
		oxygen_conc:units = "uMol L-1" ;
		oxygen_conc:valid_max = 300. ;
		oxygen_conc:valid_min = 0. ;
		oxygen_conc:_FillValue = -999. ;
	int profile_id ;
		profile_id:long_name = "Sequential Profile ID" ;
		profile_id:units = "1" ;
		profile_id:_FillValue = -127 ;
	double profile_time ;
		profile_time:long_name = "Profile Center Time" ;
		profile_time:standard_name = "time" ;
		profile_time:units = "seconds since 1970-01-01T00:00:00Z" ;
		profile_time:_FillValue = -999. ;
	double profile_lat ;
		profile_lat:long_name = "Profile Center Latitude" ;
		profile_lat:standard_name = "latitude" ;
		profile_lat:units = "degrees_north" ;
		profile_lat:_FillValue = -999. ;
	double profile_lon ;
		profile_lon:long_name = "Profile Center Longitude" ;
		profile_lon:standard_name = "longitude" ;
		profile_lon:units = "degrees_east" ;
		profile_lon:_FillValue = -999. ;

// global attributes:
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:acknowledgment = "This deployment supported the National Science Foundation and the Consortium for Ocean Leadership" ;
		:comment = "Data is not to be used for scientific purposes." ;
		:contributor_name = "John Kerfoot" ;
		:contributor_role = "Data Manager" ;
		:creator_email = "kerfoot@marine.rutgers.edu" ;
		:creator_name = "John Kerfoot" ;
		:creator_url = "http://marine.rutgers.edu/cool/auvs" ;
		:date_created = "2014-04-30T10:56:23Z" ;
		:date_issued = "2014-04-30T10:56:23Z" ;
		:date_modified = "" ;
		:format_version = "Glider_NetCDF_Profile_v1.0" ;
		:history = "/home/kerfoot/git/ooinet2epe/matlab/nc/writeOoiGliderFlatNc" ;
		:id = "" ;
		:institution = "OOI" ;
		:keywords = "AUVS > Autonomous Underwater Vehicles, Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:license = "These data were collected by the Ocean Observatory Initiative (OOI) project purely for internal system development purposes during the construction phase of the project and are offered for release to the public with no assurance of data quality, consistency, temporal continuity or additional support. The OOI Program assumes no liability resulting from the use of these data for other than the intended purpose. No data quality assurance steps have been implemented on this data to date." ;
		:metadata_link = "" ;
		:naming_authority = "edu.rutgers.marine" ;
		:platform_type = "Slocum" ;
		:processing_level = "profile" ;
		:project = "Ocean Observatories Initiative" ;
		:publisher_email = "kerfoot@marine.rutgers.edu" ;
		:publisher_name = "John Kerfoot" ;
		:publisher_url = "http://rucool.marine.rutgers.edu" ;
		:references = "http://oceanobservatories.org" ;
		:sea_name = "NE Pacific" ;
		:source = "Observational data from a profiling glider" ;
		:standard_name_vocabulary = "CF-1.6" ;
		:summary = "Observational data from an OOI Global Station Papa profiling glider" ;
		:title = "OOI GP05MOAS-GL001" ;
}
